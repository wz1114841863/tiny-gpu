`default_nettype none
`timescale 1ns/1ns

// PROGRAM COUNTER
// > Calculates the next PC for each thread to update to (but currently we assume all threads
//   update to the same PC and don't support branch divergence)
// > Currently, each thread in each core has it's own calculation for next PC
// > The NZP register value is set by the CMP instruction (based on >/=/< comparison) to
//   initiate the BRnzp instruction for branching
//   通过NZP(Negative/Zero/Positive)寄存器实现条件跳转.

/*
    1. enable: When the PC is enabled (i.e., the thread is active)
    2. core_state: When the core is in the EXECUTE state (3'b101) or UPDATE state (3'b110)
    3. decoded_nzp: The NZP bits specified in the BRnzp instruction
    4. decoded_immediate: The immediate value specified in the BRnzp instruction
    5. decoded_nzp_write_enable: When the instruction is a CMP instruction (1)
    6. decoded_pc_mux: When the instruction is a BRnzp instruction (1)
    7. alu_out: The output from the ALU used to set the NZP register
    8. current_pc: The current PC value
*/

module pc #(
    parameter DATA_MEM_DATA_BITS = 8,
    parameter PROGRAM_MEM_ADDR_BITS = 8
) (
    input wire clk,
    input wire reset,
    input wire enable, // If current block has less threads then block size, some PCs will be inactive

    // State
    input reg [2:0] core_state,

    // Control Signals
    input reg [2:0] decoded_nzp,
    input reg [DATA_MEM_DATA_BITS-1:0] decoded_immediate,
    input reg decoded_nzp_write_enable,
    input reg decoded_pc_mux,

    // ALU Output - used for alu_out[2:0] to compare with NZP register
    input reg [DATA_MEM_DATA_BITS-1:0] alu_out,

    // Current & Next PCs
    input reg [PROGRAM_MEM_ADDR_BITS-1:0] current_pc,
    output reg [PROGRAM_MEM_ADDR_BITS-1:0] next_pc
);
    reg [2:0] nzp;

    always @(posedge clk) begin
        if (reset) begin
            nzp <= 3'b0;
            next_pc <= 0;
        end else if (enable) begin
            // Update PC when core_state = EXECUTE
            if (core_state == 3'b101) begin
                if (decoded_pc_mux == 1) begin
                    if (((nzp & decoded_nzp) != 3'b0)) begin
                        // On BRnzp instruction, branch to immediate if NZP case matches previous CMP
                        next_pc <= decoded_immediate;
                    end else begin
                        // Otherwise, just update to PC + 1 (next line)
                        next_pc <= current_pc + 1;
                    end
                end else begin
                    // By default update to PC + 1 (next line)
                    next_pc <= current_pc + 1;
                end
            end

            // Store NZP when core_state = UPDATE
            // 当前NZP标志寄存器(由之前的CMP指令设置), NZP设置和分支判断之间存在一个时钟周期的延迟
            if (core_state == 3'b110) begin
                // Write to NZP register on CMP instruction
                if (decoded_nzp_write_enable) begin
                    nzp[2] <= alu_out[2];
                    nzp[1] <= alu_out[1];
                    nzp[0] <= alu_out[0];
                end
            end
        end
    end

endmodule
